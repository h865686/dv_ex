//Synchronus FIFO
